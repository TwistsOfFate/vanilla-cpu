module oz_count(
	input mode,
	input [31:0] in,
	output logic [31:0] out
);


always_comb begin
	unique case (mode)
		1'b0:
		begin
			casez (in)
				32'b00000_00000_00000_00000_00000_00000_00: out = 32'd32;
				32'b00000_00000_00000_00000_00000_00000_0?: out = 32'd31;
				32'b00000_00000_00000_00000_00000_00000_??: out = 32'd30;
				32'b00000_00000_00000_00000_00000_0000?_??: out = 32'd29;
				32'b00000_00000_00000_00000_00000_000??_??: out = 32'd28;
				32'b00000_00000_00000_00000_00000_00???_??: out = 32'd27;
				32'b00000_00000_00000_00000_00000_0????_??: out = 32'd26;
				32'b00000_00000_00000_00000_00000_?????_??: out = 32'd25;
				32'b00000_00000_00000_00000_0000?_?????_??: out = 32'd24;
				32'b00000_00000_00000_00000_000??_?????_??: out = 32'd23;
				32'b00000_00000_00000_00000_00???_?????_??: out = 32'd22;
				32'b00000_00000_00000_00000_0????_?????_??: out = 32'd21;
				32'b00000_00000_00000_00000_?????_?????_??: out = 32'd20;
				32'b00000_00000_00000_0000?_?????_?????_??: out = 32'd19;
				32'b00000_00000_00000_000??_?????_?????_??: out = 32'd18;
				32'b00000_00000_00000_00???_?????_?????_??: out = 32'd17;
				32'b00000_00000_00000_0????_?????_?????_??: out = 32'd16;
				32'b00000_00000_00000_?????_?????_?????_??: out = 32'd15;
				32'b00000_00000_0000?_?????_?????_?????_??: out = 32'd14;
				32'b00000_00000_000??_?????_?????_?????_??: out = 32'd13;
				32'b00000_00000_00???_?????_?????_?????_??: out = 32'd12;
				32'b00000_00000_0????_?????_?????_?????_??: out = 32'd11;
				32'b00000_00000_?????_?????_?????_?????_??: out = 32'd10;
				32'b00000_0000?_?????_?????_?????_?????_??: out = 32'd9;
				32'b00000_000??_?????_?????_?????_?????_??: out = 32'd8;
				32'b00000_00???_?????_?????_?????_?????_??: out = 32'd7;
				32'b00000_0????_?????_?????_?????_?????_??: out = 32'd6;
				32'b00000_?????_?????_?????_?????_?????_??: out = 32'd5;
				32'b0000?_?????_?????_?????_?????_?????_??: out = 32'd4;
				32'b000??_?????_?????_?????_?????_?????_??: out = 32'd3;
				32'b00???_?????_?????_?????_?????_?????_??: out = 32'd2;
				32'b0????_?????_?????_?????_?????_?????_??: out = 32'd1;
				default: out = 32'd0;
			endcase
		end
		1'b1:
		begin
			casez (in)
				32'b11111_11111_11111_11111_11111_11111_11: out = 32'd32;
				32'b11111_11111_11111_11111_11111_11111_1?: out = 32'd31;
				32'b11111_11111_11111_11111_11111_11111_??: out = 32'd30;
				32'b11111_11111_11111_11111_11111_1111?_??: out = 32'd29;
				32'b11111_11111_11111_11111_11111_111??_??: out = 32'd28;
				32'b11111_11111_11111_11111_11111_11???_??: out = 32'd27;
				32'b11111_11111_11111_11111_11111_1????_??: out = 32'd26;
				32'b11111_11111_11111_11111_11111_?????_??: out = 32'd25;
				32'b11111_11111_11111_11111_1111?_?????_??: out = 32'd24;
				32'b11111_11111_11111_11111_111??_?????_??: out = 32'd23;
				32'b11111_11111_11111_11111_11???_?????_??: out = 32'd22;
				32'b11111_11111_11111_11111_1????_?????_??: out = 32'd21;
				32'b11111_11111_11111_11111_?????_?????_??: out = 32'd20;
				32'b11111_11111_11111_1111?_?????_?????_??: out = 32'd19;
				32'b11111_11111_11111_111??_?????_?????_??: out = 32'd18;
				32'b11111_11111_11111_11???_?????_?????_??: out = 32'd17;
				32'b11111_11111_11111_1????_?????_?????_??: out = 32'd16;
				32'b11111_11111_11111_?????_?????_?????_??: out = 32'd15;
				32'b11111_11111_1111?_?????_?????_?????_??: out = 32'd14;
				32'b11111_11111_111??_?????_?????_?????_??: out = 32'd13;
				32'b11111_11111_11???_?????_?????_?????_??: out = 32'd12;
				32'b11111_11111_1????_?????_?????_?????_??: out = 32'd11;
				32'b11111_11111_?????_?????_?????_?????_??: out = 32'd10;
				32'b11111_1111?_?????_?????_?????_?????_??: out = 32'd9;
				32'b11111_111??_?????_?????_?????_?????_??: out = 32'd8;
				32'b11111_11???_?????_?????_?????_?????_??: out = 32'd7;
				32'b11111_1????_?????_?????_?????_?????_??: out = 32'd6;
				32'b11111_?????_?????_?????_?????_?????_??: out = 32'd5;
				32'b1111?_?????_?????_?????_?????_?????_??: out = 32'd4;
				32'b111??_?????_?????_?????_?????_?????_??: out = 32'd3;
				32'b11???_?????_?????_?????_?????_?????_??: out = 32'd2;
				32'b1????_?????_?????_?????_?????_?????_??: out = 32'd1;
				default: out = 32'd0;
			endcase
		end
	endcase
end

endmodule